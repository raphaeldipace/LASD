module InstrMemDesafio(
    input [7:0] A,
    output reg [31:0] RD
);

always @(*)
begin
    case (A)
        8'b00000000: RD = 32'b_001000_00000_00001_00000_00011_001010;
        8'b00000001: RD = 32'b_000000_00001_00001_00001_00000_100000; // *2
        8'b00000010: RD = 32'b_000000_00001_00001_00001_00000_100000; // *4
        8'b00000011: RD = 32'b_000000_00001_00001_00001_00000_100000; //*6
        8'b00000100: RD = 32'b_000000_00001_00001_00001_00000_100000; //*8
        default: RD = 32'b000000_00000_00000_00000_00000_000000; 
    endcase
end

endmodule