module mux2por1(
  input sel,
  input [7:0] a,
  input [7:0] b,
  output reg [7:0] out
);

  always @ (sel, a, b)
    case (sel)
      1'b0: out = a;
      1'b1: out = b;
      default: out = 8'hzz; // Valor indefinido padrão
    endcase
  
endmodule

